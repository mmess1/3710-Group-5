`timescale 1ns/1ps

// DE1-SoC top-level for ECE3710 ALU demo
//
// Inputs (board):
//   SW[9:0]   : use SW[7:0] as "data byte", SW[9:8] as byte select
//   KEY[0]    : reset (active-low)
//   KEY[1]    : LOAD_DATA   (active-low pulse)
//   KEY[2]    : LOAD_OPCODE (active-low pulse)
//   KEY[3]    : EXECUTE     (active-low pulse)
//
// Internal registers:
//   Rdest_reg (16), Rsrc_reg (16), Opcode_reg (8)
//   Result_reg (16), Flags_reg (5)
//
// Outputs:
//   HEX3..HEX0 : Result_reg (16-bit) as 4 hex digits
//   HEX5..HEX4 : Opcode_reg (8-bit)  as 2 hex digits
//   LEDR[4:0]  : Flags_reg [4:0]
//   LEDR[9:5]  : Opcode_reg[4:0] (quick view)

module ECE3710_top (
    input  wire        CLOCK_50,
    input  wire [9:0]  SW,
    input  wire [3:0]  KEY,
    output wire [9:0]  LEDR,
    output wire [6:0]  HEX0,
    output wire [6:0]  HEX1,
    output wire [6:0]  HEX2,
    output wire [6:0]  HEX3,
    output wire [6:0]  HEX4,
    output wire [6:0]  HEX5
);

    // Reset (KEYs are active-low)
    wire reset_n = KEY[0];

    // Button pulses (falling-edge detect on KEY1/2/3)
    wire load_data_pulse;
    wire load_op_pulse;
    wire exec_pulse;

    key_fall_pulse u_p1 (.clk(CLOCK_50), .reset_n(reset_n), .key_n(KEY[1]), .pulse(load_data_pulse));
    key_fall_pulse u_p2 (.clk(CLOCK_50), .reset_n(reset_n), .key_n(KEY[2]), .pulse(load_op_pulse));
    key_fall_pulse u_p3 (.clk(CLOCK_50), .reset_n(reset_n), .key_n(KEY[3]), .pulse(exec_pulse));

    // Input registers you "load" from switches
    reg [15:0] Rdest_reg;
    reg [15:0] Rsrc_reg;
    reg [7:0]  Opcode_reg;

    // Latched outputs for stable demo + proper WAIT/NOP behavior
    reg [15:0] Result_reg;
    reg [4:0]  Flags_reg;

    // Your ALU combinational outputs
    wire [15:0] alu_result;
    wire [4:0]  alu_flags;

    // Must match your ALU's WAIT opcode
    localparam [7:0] WAIT = 8'b0000_0000;

    // Instantiate your ALU (combinational)
    ECE3710_alu dut (
        .Rdest    (16'd2),
        .Rsrc_Imm (16'd5),
        .Opcode   (Opcode_reg),
        .Result   (alu_result),
        .Flags    (alu_flags)
    );

    // Loading/executing logic
    // SW usage:
    //   SW[7:0]  = data byte to load
    //   SW[9:8]  = which byte to load when KEY1 pressed:
    //              2'b00 -> Rdest[7:0]
    //              2'b01 -> Rdest[15:8]
    //              2'b10 -> Rsrc [7:0]
    //              2'b11 -> Rsrc [15:8]
    wire [1:0] byte_sel = SW[9:8];

    always @(posedge CLOCK_50 or negedge reset_n) begin
        if (!reset_n) begin
            Rdest_reg  <= 16'h0000;
            Rsrc_reg   <= 16'h0000;
            Opcode_reg <= 8'h00;

            Result_reg <= 16'h0000;
            Flags_reg  <= 5'b00000;
        end else begin
            // Load operand bytes
            if (load_data_pulse) begin
                case (byte_sel)
                    2'b00: Rdest_reg[7:0]   <= SW[7:0];
                    2'b01: Rdest_reg[15:8]  <= SW[7:0];
                    2'b10: Rsrc_reg[7:0]    <= SW[7:0];
                    2'b11: Rsrc_reg[15:8]   <= SW[7:0];
                    default: ;
                endcase
            end

            // Load opcode
            if (load_op_pulse) begin
                Opcode_reg <= SW[7:0];
            end

            // Execute: latch ALU outputs (WAIT/NOP holds previous)
            if (exec_pulse) begin
                if (Opcode_reg != WAIT) begin
                    Result_reg <= alu_result;
                    Flags_reg  <= alu_flags;
                end
                // else: hold Result_reg/Flags_reg
            end
        end
    end

    // LEDs: show Flags + low bits of opcode
    assign LEDR[4:0] = Flags_reg;
    //assign LEDR[9:5] = Opcode_reg[4:0];

    // 7-seg helper (active-low segments, common DE1-style)
    // If your digits appear inverted, change "assign HEXx = ..." to "~hex7(...)"
    function [6:0] hex7;
        input [3:0] x;
        begin
            case (x)
                4'h0: hex7 = 7'b1000000;
                4'h1: hex7 = 7'b1111001;
                4'h2: hex7 = 7'b0100100;
                4'h3: hex7 = 7'b0110000;
                4'h4: hex7 = 7'b0011001;
                4'h5: hex7 = 7'b0010010;
                4'h6: hex7 = 7'b0000010;
                4'h7: hex7 = 7'b1111000;
                4'h8: hex7 = 7'b0000000;
                4'h9: hex7 = 7'b0010000;
                4'hA: hex7 = 7'b0001000;
                4'hB: hex7 = 7'b0000011;
                4'hC: hex7 = 7'b1000110;
                4'hD: hex7 = 7'b0100001;
                4'hE: hex7 = 7'b0000110;
                4'hF: hex7 = 7'b0001110;
                default: hex7 = 7'b1111111;
            endcase
        end
    endfunction

    // Result on HEX3..HEX0
    assign HEX0 = hex7(Result_reg[3:0]);
    assign HEX1 = hex7(Result_reg[7:4]);
    assign HEX2 = hex7(Result_reg[11:8]);
    assign HEX3 = hex7(Result_reg[15:12]);

    // Opcode on HEX5..HEX4
    assign HEX4 = hex7(Opcode_reg[3:0]);
    assign HEX5 = hex7(Opcode_reg[7:4]);

endmodule

// Simple falling-edge pulse generator for active-low KEY buttons
// (sync + falling-edge detect; minimal debounce)
module key_fall_pulse (
    input  wire clk,
    input  wire reset_n,
    input  wire key_n,    // active-low button input
    output reg  pulse
);
    reg [2:0] sync;
    reg       prev;

    always @(posedge clk or negedge reset_n) begin
        if (!reset_n) begin
            sync  <= 3'b111;
            prev  <= 1'b1;
            pulse <= 1'b0;
        end else begin
            sync <= {sync[1:0], key_n};   // synchronize
            pulse <= (prev == 1'b1) && (sync[2] == 1'b0); // falling edge
            prev <= sync[2];
        end
    end
endmodule
